// procesador.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module procesador (
		input  wire        clk_clk,                               //                         clk.clk
		input  wire        clk_custom_in_clk,                     //               clk_custom_in.clk
		output wire        clk_custom_out_clk,                    //              clk_custom_out.clk
		output wire [31:0] divisor_clock_export,                  //               divisor_clock.export
		output wire        enable_export,                         //                      enable.export
		input  wire        fifo0_32_bit_in_valid,                 //             fifo0_32_bit_in.valid
		input  wire [31:0] fifo0_32_bit_in_data,                  //                            .data
		output wire        fifo0_32_bit_in_ready,                 //                            .ready
		input  wire        fifo0_64_bit_down_in_valid,            //        fifo0_64_bit_down_in.valid
		input  wire [31:0] fifo0_64_bit_down_in_data,             //                            .data
		output wire        fifo0_64_bit_down_in_ready,            //                            .ready
		input  wire        fifo0_64_bit_up_in_valid,              //          fifo0_64_bit_up_in.valid
		input  wire [31:0] fifo0_64_bit_up_in_data,               //                            .data
		output wire        fifo0_64_bit_up_in_ready,              //                            .ready
		input  wire        fifo1_32_bit_in_valid,                 //             fifo1_32_bit_in.valid
		input  wire [31:0] fifo1_32_bit_in_data,                  //                            .data
		output wire        fifo1_32_bit_in_ready,                 //                            .ready
		input  wire        fifo1_64_bit_down_in_valid,            //        fifo1_64_bit_down_in.valid
		input  wire [31:0] fifo1_64_bit_down_in_data,             //                            .data
		output wire        fifo1_64_bit_down_in_ready,            //                            .ready
		input  wire        fifo1_64_bit_up_in_valid,              //          fifo1_64_bit_up_in.valid
		input  wire [31:0] fifo1_64_bit_up_in_data,               //                            .data
		output wire        fifo1_64_bit_up_in_ready,              //                            .ready
		input  wire        finalizacion_export,                   //                finalizacion.export
		output wire [12:0] memory_mem_a,                          //                      memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //                            .mem_ba
		output wire        memory_mem_ck,                         //                            .mem_ck
		output wire        memory_mem_ck_n,                       //                            .mem_ck_n
		output wire        memory_mem_cke,                        //                            .mem_cke
		output wire        memory_mem_cs_n,                       //                            .mem_cs_n
		output wire        memory_mem_ras_n,                      //                            .mem_ras_n
		output wire        memory_mem_cas_n,                      //                            .mem_cas_n
		output wire        memory_mem_we_n,                       //                            .mem_we_n
		output wire        memory_mem_reset_n,                    //                            .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                         //                            .mem_dq
		inout  wire        memory_mem_dqs,                        //                            .mem_dqs
		inout  wire        memory_mem_dqs_n,                      //                            .mem_dqs_n
		output wire        memory_mem_odt,                        //                            .mem_odt
		output wire        memory_mem_dm,                         //                            .mem_dm
		input  wire        memory_oct_rzqin,                      //                            .oct_rzqin
		output wire [31:0] parameters_1_user_interface_dataout_0, // parameters_1_user_interface.dataout_0
		output wire [31:0] parameters_1_user_interface_dataout_1, //                            .dataout_1
		output wire [31:0] parameters_1_user_interface_dataout_2, //                            .dataout_2
		output wire [31:0] parameters_1_user_interface_dataout_3, //                            .dataout_3
		output wire [31:0] parameters_1_user_interface_dataout_4, //                            .dataout_4
		output wire [31:0] parameters_1_user_interface_dataout_5, //                            .dataout_5
		output wire [31:0] parameters_1_user_interface_dataout_6, //                            .dataout_6
		output wire [31:0] parameters_1_user_interface_dataout_7, //                            .dataout_7
		output wire [31:0] parameters_1_user_interface_dataout_8, //                            .dataout_8
		output wire [31:0] parameters_1_user_interface_dataout_9, //                            .dataout_9
		input  wire [31:0] parameters_1_user_interface_datain_10, //                            .datain_10
		input  wire [31:0] parameters_1_user_interface_datain_11, //                            .datain_11
		input  wire [31:0] parameters_1_user_interface_datain_12, //                            .datain_12
		input  wire [31:0] parameters_1_user_interface_datain_13, //                            .datain_13
		input  wire [31:0] parameters_1_user_interface_datain_14, //                            .datain_14
		input  wire [31:0] parameters_1_user_interface_datain_15, //                            .datain_15
		output wire [31:0] parameters_2_user_interface_dataout_0, // parameters_2_user_interface.dataout_0
		output wire [31:0] parameters_2_user_interface_dataout_1, //                            .dataout_1
		output wire [31:0] parameters_2_user_interface_dataout_2, //                            .dataout_2
		output wire [31:0] parameters_2_user_interface_dataout_3, //                            .dataout_3
		output wire [31:0] parameters_2_user_interface_dataout_4, //                            .dataout_4
		output wire [31:0] parameters_2_user_interface_dataout_5, //                            .dataout_5
		output wire [31:0] parameters_2_user_interface_dataout_6, //                            .dataout_6
		output wire [31:0] parameters_2_user_interface_dataout_7, //                            .dataout_7
		output wire [31:0] parameters_2_user_interface_dataout_8, //                            .dataout_8
		output wire [31:0] parameters_2_user_interface_dataout_9, //                            .dataout_9
		input  wire [31:0] parameters_2_user_interface_datain_10, //                            .datain_10
		input  wire [31:0] parameters_2_user_interface_datain_11, //                            .datain_11
		input  wire [31:0] parameters_2_user_interface_datain_12, //                            .datain_12
		input  wire [31:0] parameters_2_user_interface_datain_13, //                            .datain_13
		input  wire [31:0] parameters_2_user_interface_datain_14, //                            .datain_14
		input  wire [31:0] parameters_2_user_interface_datain_15, //                            .datain_15
		output wire [31:0] parameters_3_user_interface_dataout_0, // parameters_3_user_interface.dataout_0
		output wire [31:0] parameters_3_user_interface_dataout_1, //                            .dataout_1
		output wire [31:0] parameters_3_user_interface_dataout_2, //                            .dataout_2
		output wire [31:0] parameters_3_user_interface_dataout_3, //                            .dataout_3
		output wire [31:0] parameters_3_user_interface_dataout_4, //                            .dataout_4
		output wire [31:0] parameters_3_user_interface_dataout_5, //                            .dataout_5
		output wire [31:0] parameters_3_user_interface_dataout_6, //                            .dataout_6
		output wire [31:0] parameters_3_user_interface_dataout_7, //                            .dataout_7
		output wire [31:0] parameters_3_user_interface_dataout_8, //                            .dataout_8
		output wire [31:0] parameters_3_user_interface_dataout_9, //                            .dataout_9
		input  wire [31:0] parameters_3_user_interface_datain_10, //                            .datain_10
		input  wire [31:0] parameters_3_user_interface_datain_11, //                            .datain_11
		input  wire [31:0] parameters_3_user_interface_datain_12, //                            .datain_12
		input  wire [31:0] parameters_3_user_interface_datain_13, //                            .datain_13
		input  wire [31:0] parameters_3_user_interface_datain_14, //                            .datain_14
		input  wire [31:0] parameters_3_user_interface_datain_15, //                            .datain_15
		output wire [31:0] parameters_user_interface_dataout_0,   //   parameters_user_interface.dataout_0
		output wire [31:0] parameters_user_interface_dataout_1,   //                            .dataout_1
		output wire [31:0] parameters_user_interface_dataout_2,   //                            .dataout_2
		output wire [31:0] parameters_user_interface_dataout_3,   //                            .dataout_3
		output wire [31:0] parameters_user_interface_dataout_4,   //                            .dataout_4
		output wire [31:0] parameters_user_interface_dataout_5,   //                            .dataout_5
		output wire [31:0] parameters_user_interface_dataout_6,   //                            .dataout_6
		output wire [31:0] parameters_user_interface_dataout_7,   //                            .dataout_7
		output wire [31:0] parameters_user_interface_dataout_8,   //                            .dataout_8
		output wire [31:0] parameters_user_interface_dataout_9,   //                            .dataout_9
		input  wire [31:0] parameters_user_interface_datain_10,   //                            .datain_10
		input  wire [31:0] parameters_user_interface_datain_11,   //                            .datain_11
		input  wire [31:0] parameters_user_interface_datain_12,   //                            .datain_12
		input  wire [31:0] parameters_user_interface_datain_13,   //                            .datain_13
		input  wire [31:0] parameters_user_interface_datain_14,   //                            .datain_14
		input  wire [31:0] parameters_user_interface_datain_15,   //                            .datain_15
		input  wire        reset_reset_n,                         //                       reset.reset_n
		input  wire        reset_fifos_reset,                     //                 reset_fifos.reset
		output wire        reset_op_export,                       //                    reset_op.export
		input  wire [31:0] result0_32_bit_in_export,              //           result0_32_bit_in.export
		input  wire [31:0] result0_64_bit_down_in_export,         //      result0_64_bit_down_in.export
		input  wire [31:0] result0_64_bit_up_in_export,           //        result0_64_bit_up_in.export
		input  wire [31:0] result1_32_bit_in_export,              //           result1_32_bit_in.export
		input  wire [31:0] result1_64_bit_down_in_export,         //      result1_64_bit_down_in.export
		input  wire [31:0] result1_64_bit_up_in_export            //        result1_64_bit_up_in.export
	);

	wire  [63:0] pll_reconfig_from_pll_reconfig_from_pll;                          // pll:reconfig_from_pll -> pll_reconfigurar:reconfig_from_pll
	wire  [63:0] pll_reconfigurar_reconfig_to_pll_reconfig_to_pll;                 // pll_reconfigurar:reconfig_to_pll -> pll:reconfig_to_pll
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                                  // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                    // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                    // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                      // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                                   // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                    // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                      // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                                  // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                                   // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                                   // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                                   // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                                   // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                    // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                                  // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                                  // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                     // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                                   // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                                   // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                                   // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                                  // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                                   // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                                   // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                                    // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                     // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                      // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                                   // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                                  // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_readdata;    // pll_reconfigurar:mgmt_readdata -> mm_interconnect_0:pll_reconfigurar_mgmt_avalon_slave_readdata
	wire         mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_waitrequest; // pll_reconfigurar:mgmt_waitrequest -> mm_interconnect_0:pll_reconfigurar_mgmt_avalon_slave_waitrequest
	wire   [5:0] mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_address;     // mm_interconnect_0:pll_reconfigurar_mgmt_avalon_slave_address -> pll_reconfigurar:mgmt_address
	wire         mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_read;        // mm_interconnect_0:pll_reconfigurar_mgmt_avalon_slave_read -> pll_reconfigurar:mgmt_read
	wire         mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_write;       // mm_interconnect_0:pll_reconfigurar_mgmt_avalon_slave_write -> pll_reconfigurar:mgmt_write
	wire  [31:0] mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_writedata;   // mm_interconnect_0:pll_reconfigurar_mgmt_avalon_slave_writedata -> pll_reconfigurar:mgmt_writedata
	wire  [31:0] mm_interconnect_0_fifo1_32_bit_out_readdata;                      // fifo1_32_bit:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo1_32_bit_out_readdata
	wire         mm_interconnect_0_fifo1_32_bit_out_waitrequest;                   // fifo1_32_bit:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo1_32_bit_out_waitrequest
	wire   [0:0] mm_interconnect_0_fifo1_32_bit_out_address;                       // mm_interconnect_0:fifo1_32_bit_out_address -> fifo1_32_bit:avalonmm_read_slave_address
	wire         mm_interconnect_0_fifo1_32_bit_out_read;                          // mm_interconnect_0:fifo1_32_bit_out_read -> fifo1_32_bit:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo0_32_bit_out_readdata;                      // fifo0_32_bit:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo0_32_bit_out_readdata
	wire         mm_interconnect_0_fifo0_32_bit_out_waitrequest;                   // fifo0_32_bit:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo0_32_bit_out_waitrequest
	wire   [0:0] mm_interconnect_0_fifo0_32_bit_out_address;                       // mm_interconnect_0:fifo0_32_bit_out_address -> fifo0_32_bit:avalonmm_read_slave_address
	wire         mm_interconnect_0_fifo0_32_bit_out_read;                          // mm_interconnect_0:fifo0_32_bit_out_read -> fifo0_32_bit:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo1_64_bit_down_out_readdata;                 // fifo1_64_bit_down:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo1_64_bit_down_out_readdata
	wire         mm_interconnect_0_fifo1_64_bit_down_out_waitrequest;              // fifo1_64_bit_down:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo1_64_bit_down_out_waitrequest
	wire   [0:0] mm_interconnect_0_fifo1_64_bit_down_out_address;                  // mm_interconnect_0:fifo1_64_bit_down_out_address -> fifo1_64_bit_down:avalonmm_read_slave_address
	wire         mm_interconnect_0_fifo1_64_bit_down_out_read;                     // mm_interconnect_0:fifo1_64_bit_down_out_read -> fifo1_64_bit_down:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo1_64_bit_up_out_readdata;                   // fifo1_64_bit_up:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo1_64_bit_up_out_readdata
	wire         mm_interconnect_0_fifo1_64_bit_up_out_waitrequest;                // fifo1_64_bit_up:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo1_64_bit_up_out_waitrequest
	wire   [0:0] mm_interconnect_0_fifo1_64_bit_up_out_address;                    // mm_interconnect_0:fifo1_64_bit_up_out_address -> fifo1_64_bit_up:avalonmm_read_slave_address
	wire         mm_interconnect_0_fifo1_64_bit_up_out_read;                       // mm_interconnect_0:fifo1_64_bit_up_out_read -> fifo1_64_bit_up:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo0_64_bit_down_out_readdata;                 // fifo0_64_bit_down:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo0_64_bit_down_out_readdata
	wire         mm_interconnect_0_fifo0_64_bit_down_out_waitrequest;              // fifo0_64_bit_down:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo0_64_bit_down_out_waitrequest
	wire   [0:0] mm_interconnect_0_fifo0_64_bit_down_out_address;                  // mm_interconnect_0:fifo0_64_bit_down_out_address -> fifo0_64_bit_down:avalonmm_read_slave_address
	wire         mm_interconnect_0_fifo0_64_bit_down_out_read;                     // mm_interconnect_0:fifo0_64_bit_down_out_read -> fifo0_64_bit_down:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo0_64_bit_up_out_readdata;                   // fifo0_64_bit_up:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo0_64_bit_up_out_readdata
	wire         mm_interconnect_0_fifo0_64_bit_up_out_waitrequest;                // fifo0_64_bit_up:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo0_64_bit_up_out_waitrequest
	wire   [0:0] mm_interconnect_0_fifo0_64_bit_up_out_address;                    // mm_interconnect_0:fifo0_64_bit_up_out_address -> fifo0_64_bit_up:avalonmm_read_slave_address
	wire         mm_interconnect_0_fifo0_64_bit_up_out_read;                       // mm_interconnect_0:fifo0_64_bit_up_out_read -> fifo0_64_bit_up:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_parameters_3_s0_readdata;                       // parameters_3:slave_readdata -> mm_interconnect_0:parameters_3_s0_readdata
	wire   [8:0] mm_interconnect_0_parameters_3_s0_address;                        // mm_interconnect_0:parameters_3_s0_address -> parameters_3:slave_address
	wire         mm_interconnect_0_parameters_3_s0_read;                           // mm_interconnect_0:parameters_3_s0_read -> parameters_3:slave_read
	wire   [3:0] mm_interconnect_0_parameters_3_s0_byteenable;                     // mm_interconnect_0:parameters_3_s0_byteenable -> parameters_3:slave_byteenable
	wire         mm_interconnect_0_parameters_3_s0_write;                          // mm_interconnect_0:parameters_3_s0_write -> parameters_3:slave_write
	wire  [31:0] mm_interconnect_0_parameters_3_s0_writedata;                      // mm_interconnect_0:parameters_3_s0_writedata -> parameters_3:slave_writedata
	wire  [31:0] mm_interconnect_0_parameters_2_s0_readdata;                       // parameters_2:slave_readdata -> mm_interconnect_0:parameters_2_s0_readdata
	wire   [8:0] mm_interconnect_0_parameters_2_s0_address;                        // mm_interconnect_0:parameters_2_s0_address -> parameters_2:slave_address
	wire         mm_interconnect_0_parameters_2_s0_read;                           // mm_interconnect_0:parameters_2_s0_read -> parameters_2:slave_read
	wire   [3:0] mm_interconnect_0_parameters_2_s0_byteenable;                     // mm_interconnect_0:parameters_2_s0_byteenable -> parameters_2:slave_byteenable
	wire         mm_interconnect_0_parameters_2_s0_write;                          // mm_interconnect_0:parameters_2_s0_write -> parameters_2:slave_write
	wire  [31:0] mm_interconnect_0_parameters_2_s0_writedata;                      // mm_interconnect_0:parameters_2_s0_writedata -> parameters_2:slave_writedata
	wire  [31:0] mm_interconnect_0_parameters_1_s0_readdata;                       // parameters_1:slave_readdata -> mm_interconnect_0:parameters_1_s0_readdata
	wire   [8:0] mm_interconnect_0_parameters_1_s0_address;                        // mm_interconnect_0:parameters_1_s0_address -> parameters_1:slave_address
	wire         mm_interconnect_0_parameters_1_s0_read;                           // mm_interconnect_0:parameters_1_s0_read -> parameters_1:slave_read
	wire   [3:0] mm_interconnect_0_parameters_1_s0_byteenable;                     // mm_interconnect_0:parameters_1_s0_byteenable -> parameters_1:slave_byteenable
	wire         mm_interconnect_0_parameters_1_s0_write;                          // mm_interconnect_0:parameters_1_s0_write -> parameters_1:slave_write
	wire  [31:0] mm_interconnect_0_parameters_1_s0_writedata;                      // mm_interconnect_0:parameters_1_s0_writedata -> parameters_1:slave_writedata
	wire  [31:0] mm_interconnect_0_parameters_s0_readdata;                         // parameters:slave_readdata -> mm_interconnect_0:parameters_s0_readdata
	wire   [8:0] mm_interconnect_0_parameters_s0_address;                          // mm_interconnect_0:parameters_s0_address -> parameters:slave_address
	wire         mm_interconnect_0_parameters_s0_read;                             // mm_interconnect_0:parameters_s0_read -> parameters:slave_read
	wire   [3:0] mm_interconnect_0_parameters_s0_byteenable;                       // mm_interconnect_0:parameters_s0_byteenable -> parameters:slave_byteenable
	wire         mm_interconnect_0_parameters_s0_write;                            // mm_interconnect_0:parameters_s0_write -> parameters:slave_write
	wire  [31:0] mm_interconnect_0_parameters_s0_writedata;                        // mm_interconnect_0:parameters_s0_writedata -> parameters:slave_writedata
	wire  [31:0] mm_interconnect_0_result1_32_bit_s1_readdata;                     // result1_32_bit:readdata -> mm_interconnect_0:result1_32_bit_s1_readdata
	wire   [1:0] mm_interconnect_0_result1_32_bit_s1_address;                      // mm_interconnect_0:result1_32_bit_s1_address -> result1_32_bit:address
	wire  [31:0] mm_interconnect_0_result0_32_bit_s1_readdata;                     // result0_32_bit:readdata -> mm_interconnect_0:result0_32_bit_s1_readdata
	wire   [1:0] mm_interconnect_0_result0_32_bit_s1_address;                      // mm_interconnect_0:result0_32_bit_s1_address -> result0_32_bit:address
	wire  [31:0] mm_interconnect_0_result1_64_bit_down_s1_readdata;                // result1_64_bit_down:readdata -> mm_interconnect_0:result1_64_bit_down_s1_readdata
	wire   [1:0] mm_interconnect_0_result1_64_bit_down_s1_address;                 // mm_interconnect_0:result1_64_bit_down_s1_address -> result1_64_bit_down:address
	wire  [31:0] mm_interconnect_0_result1_64_bit_up_s1_readdata;                  // result1_64_bit_up:readdata -> mm_interconnect_0:result1_64_bit_up_s1_readdata
	wire   [1:0] mm_interconnect_0_result1_64_bit_up_s1_address;                   // mm_interconnect_0:result1_64_bit_up_s1_address -> result1_64_bit_up:address
	wire  [31:0] mm_interconnect_0_result0_64_bit_down_s1_readdata;                // result0_64_bit_down:readdata -> mm_interconnect_0:result0_64_bit_down_s1_readdata
	wire   [1:0] mm_interconnect_0_result0_64_bit_down_s1_address;                 // mm_interconnect_0:result0_64_bit_down_s1_address -> result0_64_bit_down:address
	wire  [31:0] mm_interconnect_0_result0_64_bit_up_s1_readdata;                  // result0_64_bit_up:readdata -> mm_interconnect_0:result0_64_bit_up_s1_readdata
	wire   [1:0] mm_interconnect_0_result0_64_bit_up_s1_address;                   // mm_interconnect_0:result0_64_bit_up_s1_address -> result0_64_bit_up:address
	wire  [31:0] mm_interconnect_0_finalizacion_s1_readdata;                       // finalizacion:readdata -> mm_interconnect_0:finalizacion_s1_readdata
	wire   [1:0] mm_interconnect_0_finalizacion_s1_address;                        // mm_interconnect_0:finalizacion_s1_address -> finalizacion:address
	wire         mm_interconnect_0_enable_s1_chipselect;                           // mm_interconnect_0:enable_s1_chipselect -> enable:chipselect
	wire  [31:0] mm_interconnect_0_enable_s1_readdata;                             // enable:readdata -> mm_interconnect_0:enable_s1_readdata
	wire   [1:0] mm_interconnect_0_enable_s1_address;                              // mm_interconnect_0:enable_s1_address -> enable:address
	wire         mm_interconnect_0_enable_s1_write;                                // mm_interconnect_0:enable_s1_write -> enable:write_n
	wire  [31:0] mm_interconnect_0_enable_s1_writedata;                            // mm_interconnect_0:enable_s1_writedata -> enable:writedata
	wire         mm_interconnect_0_reset_s1_chipselect;                            // mm_interconnect_0:reset_s1_chipselect -> reset:chipselect
	wire  [31:0] mm_interconnect_0_reset_s1_readdata;                              // reset:readdata -> mm_interconnect_0:reset_s1_readdata
	wire   [1:0] mm_interconnect_0_reset_s1_address;                               // mm_interconnect_0:reset_s1_address -> reset:address
	wire         mm_interconnect_0_reset_s1_write;                                 // mm_interconnect_0:reset_s1_write -> reset:write_n
	wire  [31:0] mm_interconnect_0_reset_s1_writedata;                             // mm_interconnect_0:reset_s1_writedata -> reset:writedata
	wire         mm_interconnect_0_divisor_clock_s1_chipselect;                    // mm_interconnect_0:divisor_clock_s1_chipselect -> divisor_clock:chipselect
	wire  [31:0] mm_interconnect_0_divisor_clock_s1_readdata;                      // divisor_clock:readdata -> mm_interconnect_0:divisor_clock_s1_readdata
	wire   [1:0] mm_interconnect_0_divisor_clock_s1_address;                       // mm_interconnect_0:divisor_clock_s1_address -> divisor_clock:address
	wire         mm_interconnect_0_divisor_clock_s1_write;                         // mm_interconnect_0:divisor_clock_s1_write -> divisor_clock:write_n
	wire  [31:0] mm_interconnect_0_divisor_clock_s1_writedata;                     // mm_interconnect_0:divisor_clock_s1_writedata -> divisor_clock:writedata
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [divisor_clock:reset_n, enable:reset_n, finalizacion:reset_n, mm_interconnect_0:pll_reconfigurar_mgmt_reset_reset_bridge_in_reset_reset, parameters:reset, parameters_1:reset, parameters_2:reset, parameters_3:reset, pll_reconfigurar:mgmt_reset, result0_32_bit:reset_n, result0_64_bit_down:reset_n, result0_64_bit_up:reset_n, result1_32_bit:reset_n, result1_64_bit_down:reset_n, result1_64_bit_up:reset_n]
	wire         rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> [fifo0_32_bit:reset_n, fifo0_64_bit_down:reset_n, fifo0_64_bit_up:reset_n, fifo1_32_bit:reset_n, fifo1_64_bit_down:reset_n, fifo1_64_bit_up:reset_n, mm_interconnect_0:fifo1_32_bit_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                               // rst_controller_002:reset_out -> [mm_interconnect_0:reset_reset_reset_bridge_in_reset_reset, reset:reset_n]
	wire         rst_controller_003_reset_out_reset;                               // rst_controller_003:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                                            // hps_0:h2f_rst_n -> rst_controller_003:reset_in0

	procesador_divisor_clock divisor_clock (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_divisor_clock_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_divisor_clock_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_divisor_clock_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_divisor_clock_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_divisor_clock_s1_readdata),   //                    .readdata
		.out_port   (divisor_clock_export)                           // external_connection.export
	);

	procesador_enable enable (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_enable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_enable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_enable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_enable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_enable_s1_readdata),   //                    .readdata
		.out_port   (enable_export)                           // external_connection.export
	);

	procesador_fifo0_32_bit fifo0_32_bit (
		.wrclock                         (clk_custom_in_clk),                              //   clk_in.clk
		.reset_n                         (~rst_controller_001_reset_out_reset),            // reset_in.reset_n
		.avalonst_sink_valid             (fifo0_32_bit_in_valid),                          //       in.valid
		.avalonst_sink_data              (fifo0_32_bit_in_data),                           //         .data
		.avalonst_sink_ready             (fifo0_32_bit_in_ready),                          //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_fifo0_32_bit_out_readdata),    //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_fifo0_32_bit_out_read),        //         .read
		.avalonmm_read_slave_address     (mm_interconnect_0_fifo0_32_bit_out_address),     //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_fifo0_32_bit_out_waitrequest)  //         .waitrequest
	);

	procesador_fifo0_64_bit_down fifo0_64_bit_down (
		.wrclock                         (clk_custom_in_clk),                                   //   clk_in.clk
		.reset_n                         (~rst_controller_001_reset_out_reset),                 // reset_in.reset_n
		.avalonst_sink_valid             (fifo0_64_bit_down_in_valid),                          //       in.valid
		.avalonst_sink_data              (fifo0_64_bit_down_in_data),                           //         .data
		.avalonst_sink_ready             (fifo0_64_bit_down_in_ready),                          //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_fifo0_64_bit_down_out_readdata),    //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_fifo0_64_bit_down_out_read),        //         .read
		.avalonmm_read_slave_address     (mm_interconnect_0_fifo0_64_bit_down_out_address),     //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_fifo0_64_bit_down_out_waitrequest)  //         .waitrequest
	);

	procesador_fifo0_64_bit_down fifo0_64_bit_up (
		.wrclock                         (clk_custom_in_clk),                                 //   clk_in.clk
		.reset_n                         (~rst_controller_001_reset_out_reset),               // reset_in.reset_n
		.avalonst_sink_valid             (fifo0_64_bit_up_in_valid),                          //       in.valid
		.avalonst_sink_data              (fifo0_64_bit_up_in_data),                           //         .data
		.avalonst_sink_ready             (fifo0_64_bit_up_in_ready),                          //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_fifo0_64_bit_up_out_readdata),    //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_fifo0_64_bit_up_out_read),        //         .read
		.avalonmm_read_slave_address     (mm_interconnect_0_fifo0_64_bit_up_out_address),     //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_fifo0_64_bit_up_out_waitrequest)  //         .waitrequest
	);

	procesador_fifo0_32_bit fifo1_32_bit (
		.wrclock                         (clk_custom_in_clk),                              //   clk_in.clk
		.reset_n                         (~rst_controller_001_reset_out_reset),            // reset_in.reset_n
		.avalonst_sink_valid             (fifo1_32_bit_in_valid),                          //       in.valid
		.avalonst_sink_data              (fifo1_32_bit_in_data),                           //         .data
		.avalonst_sink_ready             (fifo1_32_bit_in_ready),                          //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_fifo1_32_bit_out_readdata),    //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_fifo1_32_bit_out_read),        //         .read
		.avalonmm_read_slave_address     (mm_interconnect_0_fifo1_32_bit_out_address),     //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_fifo1_32_bit_out_waitrequest)  //         .waitrequest
	);

	procesador_fifo0_64_bit_down fifo1_64_bit_down (
		.wrclock                         (clk_custom_in_clk),                                   //   clk_in.clk
		.reset_n                         (~rst_controller_001_reset_out_reset),                 // reset_in.reset_n
		.avalonst_sink_valid             (fifo1_64_bit_down_in_valid),                          //       in.valid
		.avalonst_sink_data              (fifo1_64_bit_down_in_data),                           //         .data
		.avalonst_sink_ready             (fifo1_64_bit_down_in_ready),                          //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_fifo1_64_bit_down_out_readdata),    //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_fifo1_64_bit_down_out_read),        //         .read
		.avalonmm_read_slave_address     (mm_interconnect_0_fifo1_64_bit_down_out_address),     //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_fifo1_64_bit_down_out_waitrequest)  //         .waitrequest
	);

	procesador_fifo0_64_bit_down fifo1_64_bit_up (
		.wrclock                         (clk_custom_in_clk),                                 //   clk_in.clk
		.reset_n                         (~rst_controller_001_reset_out_reset),               // reset_in.reset_n
		.avalonst_sink_valid             (fifo1_64_bit_up_in_valid),                          //       in.valid
		.avalonst_sink_data              (fifo1_64_bit_up_in_data),                           //         .data
		.avalonst_sink_ready             (fifo1_64_bit_up_in_ready),                          //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_fifo1_64_bit_up_out_readdata),    //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_fifo1_64_bit_up_out_read),        //         .read
		.avalonmm_read_slave_address     (mm_interconnect_0_fifo1_64_bit_up_out_address),     //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_fifo1_64_bit_up_out_waitrequest)  //         .waitrequest
	);

	procesador_finalizacion finalizacion (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_finalizacion_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_finalizacion_s1_readdata), //                    .readdata
		.in_port  (finalizacion_export)                         // external_connection.export
	);

	procesador_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.mem_a          (memory_mem_a),                    //            memory.mem_a
		.mem_ba         (memory_mem_ba),                   //                  .mem_ba
		.mem_ck         (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n       (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke        (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n       (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n      (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n      (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n       (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n    (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq         (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs        (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n      (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt        (memory_mem_odt),                  //                  .mem_odt
		.mem_dm         (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin      (memory_oct_rzqin),                //                  .oct_rzqin
		.h2f_rst_n      (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_lw_axi_clk (clk_clk),                         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID    (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR  (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN   (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE  (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK  (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT  (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID     (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA   (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB   (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST   (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID  (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY  (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID     (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP   (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID  (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY  (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID    (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR  (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN   (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE  (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK  (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT  (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID     (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA   (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP   (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST   (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID  (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY  (hps_0_h2f_lw_axi_master_rready)   //                  .rready
	);

	slave_template #(
		.DATA_WIDTH          (32),
		.ENABLE_SYNC_SIGNALS (0),
		.MODE_0              (0),
		.MODE_1              (0),
		.MODE_2              (0),
		.MODE_3              (0),
		.MODE_4              (0),
		.MODE_5              (0),
		.MODE_6              (0),
		.MODE_7              (0),
		.MODE_8              (0),
		.MODE_9              (0),
		.MODE_10             (1),
		.MODE_11             (1),
		.MODE_12             (1),
		.MODE_13             (1),
		.MODE_14             (1),
		.MODE_15             (1),
		.IRQ_EN              (0)
	) parameters (
		.clk              (clk_clk),                                    //       clock_reset.clk
		.reset            (rst_controller_reset_out_reset),             // clock_reset_reset.reset
		.slave_address    (mm_interconnect_0_parameters_s0_address),    //                s0.address
		.slave_read       (mm_interconnect_0_parameters_s0_read),       //                  .read
		.slave_write      (mm_interconnect_0_parameters_s0_write),      //                  .write
		.slave_readdata   (mm_interconnect_0_parameters_s0_readdata),   //                  .readdata
		.slave_writedata  (mm_interconnect_0_parameters_s0_writedata),  //                  .writedata
		.slave_byteenable (mm_interconnect_0_parameters_s0_byteenable), //                  .byteenable
		.user_dataout_0   (parameters_user_interface_dataout_0),        //    user_interface.export
		.user_dataout_1   (parameters_user_interface_dataout_1),        //                  .export
		.user_dataout_2   (parameters_user_interface_dataout_2),        //                  .export
		.user_dataout_3   (parameters_user_interface_dataout_3),        //                  .export
		.user_dataout_4   (parameters_user_interface_dataout_4),        //                  .export
		.user_dataout_5   (parameters_user_interface_dataout_5),        //                  .export
		.user_dataout_6   (parameters_user_interface_dataout_6),        //                  .export
		.user_dataout_7   (parameters_user_interface_dataout_7),        //                  .export
		.user_dataout_8   (parameters_user_interface_dataout_8),        //                  .export
		.user_dataout_9   (parameters_user_interface_dataout_9),        //                  .export
		.user_datain_10   (parameters_user_interface_datain_10),        //                  .export
		.user_datain_11   (parameters_user_interface_datain_11),        //                  .export
		.user_datain_12   (parameters_user_interface_datain_12),        //                  .export
		.user_datain_13   (parameters_user_interface_datain_13),        //                  .export
		.user_datain_14   (parameters_user_interface_datain_14),        //                  .export
		.user_datain_15   (parameters_user_interface_datain_15),        //                  .export
		.slave_irq        (),                                           //       (terminated)
		.user_dataout_10  (),                                           //       (terminated)
		.user_dataout_11  (),                                           //       (terminated)
		.user_dataout_12  (),                                           //       (terminated)
		.user_dataout_13  (),                                           //       (terminated)
		.user_dataout_14  (),                                           //       (terminated)
		.user_dataout_15  (),                                           //       (terminated)
		.user_datain_0    (32'b00000000000000000000000000000000),       //       (terminated)
		.user_datain_1    (32'b00000000000000000000000000000000),       //       (terminated)
		.user_datain_2    (32'b00000000000000000000000000000000),       //       (terminated)
		.user_datain_3    (32'b00000000000000000000000000000000),       //       (terminated)
		.user_datain_4    (32'b00000000000000000000000000000000),       //       (terminated)
		.user_datain_5    (32'b00000000000000000000000000000000),       //       (terminated)
		.user_datain_6    (32'b00000000000000000000000000000000),       //       (terminated)
		.user_datain_7    (32'b00000000000000000000000000000000),       //       (terminated)
		.user_datain_8    (32'b00000000000000000000000000000000),       //       (terminated)
		.user_datain_9    (32'b00000000000000000000000000000000),       //       (terminated)
		.user_write       (),                                           //       (terminated)
		.user_read        (),                                           //       (terminated)
		.user_chipselect  ()                                            //       (terminated)
	);

	slave_template #(
		.DATA_WIDTH          (32),
		.ENABLE_SYNC_SIGNALS (0),
		.MODE_0              (0),
		.MODE_1              (0),
		.MODE_2              (0),
		.MODE_3              (0),
		.MODE_4              (0),
		.MODE_5              (0),
		.MODE_6              (0),
		.MODE_7              (0),
		.MODE_8              (0),
		.MODE_9              (0),
		.MODE_10             (1),
		.MODE_11             (1),
		.MODE_12             (1),
		.MODE_13             (1),
		.MODE_14             (1),
		.MODE_15             (1),
		.IRQ_EN              (0)
	) parameters_1 (
		.clk              (clk_clk),                                      //       clock_reset.clk
		.reset            (rst_controller_reset_out_reset),               // clock_reset_reset.reset
		.slave_address    (mm_interconnect_0_parameters_1_s0_address),    //                s0.address
		.slave_read       (mm_interconnect_0_parameters_1_s0_read),       //                  .read
		.slave_write      (mm_interconnect_0_parameters_1_s0_write),      //                  .write
		.slave_readdata   (mm_interconnect_0_parameters_1_s0_readdata),   //                  .readdata
		.slave_writedata  (mm_interconnect_0_parameters_1_s0_writedata),  //                  .writedata
		.slave_byteenable (mm_interconnect_0_parameters_1_s0_byteenable), //                  .byteenable
		.user_dataout_0   (parameters_1_user_interface_dataout_0),        //    user_interface.export
		.user_dataout_1   (parameters_1_user_interface_dataout_1),        //                  .export
		.user_dataout_2   (parameters_1_user_interface_dataout_2),        //                  .export
		.user_dataout_3   (parameters_1_user_interface_dataout_3),        //                  .export
		.user_dataout_4   (parameters_1_user_interface_dataout_4),        //                  .export
		.user_dataout_5   (parameters_1_user_interface_dataout_5),        //                  .export
		.user_dataout_6   (parameters_1_user_interface_dataout_6),        //                  .export
		.user_dataout_7   (parameters_1_user_interface_dataout_7),        //                  .export
		.user_dataout_8   (parameters_1_user_interface_dataout_8),        //                  .export
		.user_dataout_9   (parameters_1_user_interface_dataout_9),        //                  .export
		.user_datain_10   (parameters_1_user_interface_datain_10),        //                  .export
		.user_datain_11   (parameters_1_user_interface_datain_11),        //                  .export
		.user_datain_12   (parameters_1_user_interface_datain_12),        //                  .export
		.user_datain_13   (parameters_1_user_interface_datain_13),        //                  .export
		.user_datain_14   (parameters_1_user_interface_datain_14),        //                  .export
		.user_datain_15   (parameters_1_user_interface_datain_15),        //                  .export
		.slave_irq        (),                                             //       (terminated)
		.user_dataout_10  (),                                             //       (terminated)
		.user_dataout_11  (),                                             //       (terminated)
		.user_dataout_12  (),                                             //       (terminated)
		.user_dataout_13  (),                                             //       (terminated)
		.user_dataout_14  (),                                             //       (terminated)
		.user_dataout_15  (),                                             //       (terminated)
		.user_datain_0    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_1    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_2    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_3    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_4    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_5    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_6    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_7    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_8    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_9    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_write       (),                                             //       (terminated)
		.user_read        (),                                             //       (terminated)
		.user_chipselect  ()                                              //       (terminated)
	);

	slave_template #(
		.DATA_WIDTH          (32),
		.ENABLE_SYNC_SIGNALS (0),
		.MODE_0              (0),
		.MODE_1              (0),
		.MODE_2              (0),
		.MODE_3              (0),
		.MODE_4              (0),
		.MODE_5              (0),
		.MODE_6              (0),
		.MODE_7              (0),
		.MODE_8              (0),
		.MODE_9              (0),
		.MODE_10             (1),
		.MODE_11             (1),
		.MODE_12             (1),
		.MODE_13             (1),
		.MODE_14             (1),
		.MODE_15             (1),
		.IRQ_EN              (0)
	) parameters_2 (
		.clk              (clk_clk),                                      //       clock_reset.clk
		.reset            (rst_controller_reset_out_reset),               // clock_reset_reset.reset
		.slave_address    (mm_interconnect_0_parameters_2_s0_address),    //                s0.address
		.slave_read       (mm_interconnect_0_parameters_2_s0_read),       //                  .read
		.slave_write      (mm_interconnect_0_parameters_2_s0_write),      //                  .write
		.slave_readdata   (mm_interconnect_0_parameters_2_s0_readdata),   //                  .readdata
		.slave_writedata  (mm_interconnect_0_parameters_2_s0_writedata),  //                  .writedata
		.slave_byteenable (mm_interconnect_0_parameters_2_s0_byteenable), //                  .byteenable
		.user_dataout_0   (parameters_2_user_interface_dataout_0),        //    user_interface.export
		.user_dataout_1   (parameters_2_user_interface_dataout_1),        //                  .export
		.user_dataout_2   (parameters_2_user_interface_dataout_2),        //                  .export
		.user_dataout_3   (parameters_2_user_interface_dataout_3),        //                  .export
		.user_dataout_4   (parameters_2_user_interface_dataout_4),        //                  .export
		.user_dataout_5   (parameters_2_user_interface_dataout_5),        //                  .export
		.user_dataout_6   (parameters_2_user_interface_dataout_6),        //                  .export
		.user_dataout_7   (parameters_2_user_interface_dataout_7),        //                  .export
		.user_dataout_8   (parameters_2_user_interface_dataout_8),        //                  .export
		.user_dataout_9   (parameters_2_user_interface_dataout_9),        //                  .export
		.user_datain_10   (parameters_2_user_interface_datain_10),        //                  .export
		.user_datain_11   (parameters_2_user_interface_datain_11),        //                  .export
		.user_datain_12   (parameters_2_user_interface_datain_12),        //                  .export
		.user_datain_13   (parameters_2_user_interface_datain_13),        //                  .export
		.user_datain_14   (parameters_2_user_interface_datain_14),        //                  .export
		.user_datain_15   (parameters_2_user_interface_datain_15),        //                  .export
		.slave_irq        (),                                             //       (terminated)
		.user_dataout_10  (),                                             //       (terminated)
		.user_dataout_11  (),                                             //       (terminated)
		.user_dataout_12  (),                                             //       (terminated)
		.user_dataout_13  (),                                             //       (terminated)
		.user_dataout_14  (),                                             //       (terminated)
		.user_dataout_15  (),                                             //       (terminated)
		.user_datain_0    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_1    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_2    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_3    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_4    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_5    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_6    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_7    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_8    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_9    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_write       (),                                             //       (terminated)
		.user_read        (),                                             //       (terminated)
		.user_chipselect  ()                                              //       (terminated)
	);

	slave_template #(
		.DATA_WIDTH          (32),
		.ENABLE_SYNC_SIGNALS (0),
		.MODE_0              (0),
		.MODE_1              (0),
		.MODE_2              (0),
		.MODE_3              (0),
		.MODE_4              (0),
		.MODE_5              (0),
		.MODE_6              (0),
		.MODE_7              (0),
		.MODE_8              (0),
		.MODE_9              (0),
		.MODE_10             (1),
		.MODE_11             (1),
		.MODE_12             (1),
		.MODE_13             (1),
		.MODE_14             (1),
		.MODE_15             (1),
		.IRQ_EN              (0)
	) parameters_3 (
		.clk              (clk_clk),                                      //       clock_reset.clk
		.reset            (rst_controller_reset_out_reset),               // clock_reset_reset.reset
		.slave_address    (mm_interconnect_0_parameters_3_s0_address),    //                s0.address
		.slave_read       (mm_interconnect_0_parameters_3_s0_read),       //                  .read
		.slave_write      (mm_interconnect_0_parameters_3_s0_write),      //                  .write
		.slave_readdata   (mm_interconnect_0_parameters_3_s0_readdata),   //                  .readdata
		.slave_writedata  (mm_interconnect_0_parameters_3_s0_writedata),  //                  .writedata
		.slave_byteenable (mm_interconnect_0_parameters_3_s0_byteenable), //                  .byteenable
		.user_dataout_0   (parameters_3_user_interface_dataout_0),        //    user_interface.export
		.user_dataout_1   (parameters_3_user_interface_dataout_1),        //                  .export
		.user_dataout_2   (parameters_3_user_interface_dataout_2),        //                  .export
		.user_dataout_3   (parameters_3_user_interface_dataout_3),        //                  .export
		.user_dataout_4   (parameters_3_user_interface_dataout_4),        //                  .export
		.user_dataout_5   (parameters_3_user_interface_dataout_5),        //                  .export
		.user_dataout_6   (parameters_3_user_interface_dataout_6),        //                  .export
		.user_dataout_7   (parameters_3_user_interface_dataout_7),        //                  .export
		.user_dataout_8   (parameters_3_user_interface_dataout_8),        //                  .export
		.user_dataout_9   (parameters_3_user_interface_dataout_9),        //                  .export
		.user_datain_10   (parameters_3_user_interface_datain_10),        //                  .export
		.user_datain_11   (parameters_3_user_interface_datain_11),        //                  .export
		.user_datain_12   (parameters_3_user_interface_datain_12),        //                  .export
		.user_datain_13   (parameters_3_user_interface_datain_13),        //                  .export
		.user_datain_14   (parameters_3_user_interface_datain_14),        //                  .export
		.user_datain_15   (parameters_3_user_interface_datain_15),        //                  .export
		.slave_irq        (),                                             //       (terminated)
		.user_dataout_10  (),                                             //       (terminated)
		.user_dataout_11  (),                                             //       (terminated)
		.user_dataout_12  (),                                             //       (terminated)
		.user_dataout_13  (),                                             //       (terminated)
		.user_dataout_14  (),                                             //       (terminated)
		.user_dataout_15  (),                                             //       (terminated)
		.user_datain_0    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_1    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_2    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_3    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_4    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_5    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_6    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_7    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_8    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_datain_9    (32'b00000000000000000000000000000000),         //       (terminated)
		.user_write       (),                                             //       (terminated)
		.user_read        (),                                             //       (terminated)
		.user_chipselect  ()                                              //       (terminated)
	);

	procesador_pll pll (
		.refclk            (clk_clk),                                          //            refclk.clk
		.rst               (~reset_reset_n),                                   //             reset.reset
		.outclk_0          (clk_custom_out_clk),                               //           outclk0.clk
		.reconfig_to_pll   (pll_reconfigurar_reconfig_to_pll_reconfig_to_pll), //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_reconfig_from_pll_reconfig_from_pll),          // reconfig_from_pll.reconfig_from_pll
		.locked            ()                                                  //       (terminated)
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_reconfigurar (
		.mgmt_clk          (clk_clk),                                                          //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_reset_out_reset),                                   //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pll_reconfigurar_reconfig_to_pll_reconfig_to_pll),                 //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_reconfig_from_pll_reconfig_from_pll),                          // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                           //       (terminated)
	);

	procesador_reset reset (
		.clk        (clk_custom_in_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reset_s1_readdata),   //                    .readdata
		.out_port   (reset_op_export)                        // external_connection.export
	);

	procesador_result0_32_bit result0_32_bit (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_result0_32_bit_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_result0_32_bit_s1_readdata), //                    .readdata
		.in_port  (result0_32_bit_in_export)                      // external_connection.export
	);

	procesador_result0_32_bit result0_64_bit_down (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (mm_interconnect_0_result0_64_bit_down_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_result0_64_bit_down_s1_readdata), //                    .readdata
		.in_port  (result0_64_bit_down_in_export)                      // external_connection.export
	);

	procesador_result0_32_bit result0_64_bit_up (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_result0_64_bit_up_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_result0_64_bit_up_s1_readdata), //                    .readdata
		.in_port  (result0_64_bit_up_in_export)                      // external_connection.export
	);

	procesador_result0_32_bit result1_32_bit (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_result1_32_bit_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_result1_32_bit_s1_readdata), //                    .readdata
		.in_port  (result1_32_bit_in_export)                      // external_connection.export
	);

	procesador_result0_32_bit result1_64_bit_down (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (mm_interconnect_0_result1_64_bit_down_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_result1_64_bit_down_s1_readdata), //                    .readdata
		.in_port  (result1_64_bit_down_in_export)                      // external_connection.export
	);

	procesador_result0_32_bit result1_64_bit_up (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_result1_64_bit_up_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_result1_64_bit_up_s1_readdata), //                    .readdata
		.in_port  (result1_64_bit_up_in_export)                      // external_connection.export
	);

	procesador_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                     //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                                   //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                                    //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                                   //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                                  //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                                   //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                                  //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                                   //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                                  //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                                  //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                      //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                                    //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                                    //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                                    //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                                   //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                                   //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                      //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                                    //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                                   //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                                   //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                     //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                                   //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                                    //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                                   //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                                  //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                                   //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                                  //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                                   //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                                  //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                                  //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                      //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                                    //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                                    //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                                    //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                                   //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                                   //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                          //                                                     clk_0_clk.clk
		.clock_bridge_0_out_clk_clk                                          (clk_custom_in_clk),                                                //                                        clock_bridge_0_out_clk.clk
		.fifo1_32_bit_reset_in_reset_bridge_in_reset_reset                   (rst_controller_001_reset_out_reset),                               //                   fifo1_32_bit_reset_in_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                               // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.pll_reconfigurar_mgmt_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                   //             pll_reconfigurar_mgmt_reset_reset_bridge_in_reset.reset
		.reset_reset_reset_bridge_in_reset_reset                             (rst_controller_002_reset_out_reset),                               //                             reset_reset_reset_bridge_in_reset.reset
		.divisor_clock_s1_address                                            (mm_interconnect_0_divisor_clock_s1_address),                       //                                              divisor_clock_s1.address
		.divisor_clock_s1_write                                              (mm_interconnect_0_divisor_clock_s1_write),                         //                                                              .write
		.divisor_clock_s1_readdata                                           (mm_interconnect_0_divisor_clock_s1_readdata),                      //                                                              .readdata
		.divisor_clock_s1_writedata                                          (mm_interconnect_0_divisor_clock_s1_writedata),                     //                                                              .writedata
		.divisor_clock_s1_chipselect                                         (mm_interconnect_0_divisor_clock_s1_chipselect),                    //                                                              .chipselect
		.enable_s1_address                                                   (mm_interconnect_0_enable_s1_address),                              //                                                     enable_s1.address
		.enable_s1_write                                                     (mm_interconnect_0_enable_s1_write),                                //                                                              .write
		.enable_s1_readdata                                                  (mm_interconnect_0_enable_s1_readdata),                             //                                                              .readdata
		.enable_s1_writedata                                                 (mm_interconnect_0_enable_s1_writedata),                            //                                                              .writedata
		.enable_s1_chipselect                                                (mm_interconnect_0_enable_s1_chipselect),                           //                                                              .chipselect
		.fifo0_32_bit_out_address                                            (mm_interconnect_0_fifo0_32_bit_out_address),                       //                                              fifo0_32_bit_out.address
		.fifo0_32_bit_out_read                                               (mm_interconnect_0_fifo0_32_bit_out_read),                          //                                                              .read
		.fifo0_32_bit_out_readdata                                           (mm_interconnect_0_fifo0_32_bit_out_readdata),                      //                                                              .readdata
		.fifo0_32_bit_out_waitrequest                                        (mm_interconnect_0_fifo0_32_bit_out_waitrequest),                   //                                                              .waitrequest
		.fifo0_64_bit_down_out_address                                       (mm_interconnect_0_fifo0_64_bit_down_out_address),                  //                                         fifo0_64_bit_down_out.address
		.fifo0_64_bit_down_out_read                                          (mm_interconnect_0_fifo0_64_bit_down_out_read),                     //                                                              .read
		.fifo0_64_bit_down_out_readdata                                      (mm_interconnect_0_fifo0_64_bit_down_out_readdata),                 //                                                              .readdata
		.fifo0_64_bit_down_out_waitrequest                                   (mm_interconnect_0_fifo0_64_bit_down_out_waitrequest),              //                                                              .waitrequest
		.fifo0_64_bit_up_out_address                                         (mm_interconnect_0_fifo0_64_bit_up_out_address),                    //                                           fifo0_64_bit_up_out.address
		.fifo0_64_bit_up_out_read                                            (mm_interconnect_0_fifo0_64_bit_up_out_read),                       //                                                              .read
		.fifo0_64_bit_up_out_readdata                                        (mm_interconnect_0_fifo0_64_bit_up_out_readdata),                   //                                                              .readdata
		.fifo0_64_bit_up_out_waitrequest                                     (mm_interconnect_0_fifo0_64_bit_up_out_waitrequest),                //                                                              .waitrequest
		.fifo1_32_bit_out_address                                            (mm_interconnect_0_fifo1_32_bit_out_address),                       //                                              fifo1_32_bit_out.address
		.fifo1_32_bit_out_read                                               (mm_interconnect_0_fifo1_32_bit_out_read),                          //                                                              .read
		.fifo1_32_bit_out_readdata                                           (mm_interconnect_0_fifo1_32_bit_out_readdata),                      //                                                              .readdata
		.fifo1_32_bit_out_waitrequest                                        (mm_interconnect_0_fifo1_32_bit_out_waitrequest),                   //                                                              .waitrequest
		.fifo1_64_bit_down_out_address                                       (mm_interconnect_0_fifo1_64_bit_down_out_address),                  //                                         fifo1_64_bit_down_out.address
		.fifo1_64_bit_down_out_read                                          (mm_interconnect_0_fifo1_64_bit_down_out_read),                     //                                                              .read
		.fifo1_64_bit_down_out_readdata                                      (mm_interconnect_0_fifo1_64_bit_down_out_readdata),                 //                                                              .readdata
		.fifo1_64_bit_down_out_waitrequest                                   (mm_interconnect_0_fifo1_64_bit_down_out_waitrequest),              //                                                              .waitrequest
		.fifo1_64_bit_up_out_address                                         (mm_interconnect_0_fifo1_64_bit_up_out_address),                    //                                           fifo1_64_bit_up_out.address
		.fifo1_64_bit_up_out_read                                            (mm_interconnect_0_fifo1_64_bit_up_out_read),                       //                                                              .read
		.fifo1_64_bit_up_out_readdata                                        (mm_interconnect_0_fifo1_64_bit_up_out_readdata),                   //                                                              .readdata
		.fifo1_64_bit_up_out_waitrequest                                     (mm_interconnect_0_fifo1_64_bit_up_out_waitrequest),                //                                                              .waitrequest
		.finalizacion_s1_address                                             (mm_interconnect_0_finalizacion_s1_address),                        //                                               finalizacion_s1.address
		.finalizacion_s1_readdata                                            (mm_interconnect_0_finalizacion_s1_readdata),                       //                                                              .readdata
		.parameters_s0_address                                               (mm_interconnect_0_parameters_s0_address),                          //                                                 parameters_s0.address
		.parameters_s0_write                                                 (mm_interconnect_0_parameters_s0_write),                            //                                                              .write
		.parameters_s0_read                                                  (mm_interconnect_0_parameters_s0_read),                             //                                                              .read
		.parameters_s0_readdata                                              (mm_interconnect_0_parameters_s0_readdata),                         //                                                              .readdata
		.parameters_s0_writedata                                             (mm_interconnect_0_parameters_s0_writedata),                        //                                                              .writedata
		.parameters_s0_byteenable                                            (mm_interconnect_0_parameters_s0_byteenable),                       //                                                              .byteenable
		.parameters_1_s0_address                                             (mm_interconnect_0_parameters_1_s0_address),                        //                                               parameters_1_s0.address
		.parameters_1_s0_write                                               (mm_interconnect_0_parameters_1_s0_write),                          //                                                              .write
		.parameters_1_s0_read                                                (mm_interconnect_0_parameters_1_s0_read),                           //                                                              .read
		.parameters_1_s0_readdata                                            (mm_interconnect_0_parameters_1_s0_readdata),                       //                                                              .readdata
		.parameters_1_s0_writedata                                           (mm_interconnect_0_parameters_1_s0_writedata),                      //                                                              .writedata
		.parameters_1_s0_byteenable                                          (mm_interconnect_0_parameters_1_s0_byteenable),                     //                                                              .byteenable
		.parameters_2_s0_address                                             (mm_interconnect_0_parameters_2_s0_address),                        //                                               parameters_2_s0.address
		.parameters_2_s0_write                                               (mm_interconnect_0_parameters_2_s0_write),                          //                                                              .write
		.parameters_2_s0_read                                                (mm_interconnect_0_parameters_2_s0_read),                           //                                                              .read
		.parameters_2_s0_readdata                                            (mm_interconnect_0_parameters_2_s0_readdata),                       //                                                              .readdata
		.parameters_2_s0_writedata                                           (mm_interconnect_0_parameters_2_s0_writedata),                      //                                                              .writedata
		.parameters_2_s0_byteenable                                          (mm_interconnect_0_parameters_2_s0_byteenable),                     //                                                              .byteenable
		.parameters_3_s0_address                                             (mm_interconnect_0_parameters_3_s0_address),                        //                                               parameters_3_s0.address
		.parameters_3_s0_write                                               (mm_interconnect_0_parameters_3_s0_write),                          //                                                              .write
		.parameters_3_s0_read                                                (mm_interconnect_0_parameters_3_s0_read),                           //                                                              .read
		.parameters_3_s0_readdata                                            (mm_interconnect_0_parameters_3_s0_readdata),                       //                                                              .readdata
		.parameters_3_s0_writedata                                           (mm_interconnect_0_parameters_3_s0_writedata),                      //                                                              .writedata
		.parameters_3_s0_byteenable                                          (mm_interconnect_0_parameters_3_s0_byteenable),                     //                                                              .byteenable
		.pll_reconfigurar_mgmt_avalon_slave_address                          (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_address),     //                            pll_reconfigurar_mgmt_avalon_slave.address
		.pll_reconfigurar_mgmt_avalon_slave_write                            (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_write),       //                                                              .write
		.pll_reconfigurar_mgmt_avalon_slave_read                             (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_read),        //                                                              .read
		.pll_reconfigurar_mgmt_avalon_slave_readdata                         (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_readdata),    //                                                              .readdata
		.pll_reconfigurar_mgmt_avalon_slave_writedata                        (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_writedata),   //                                                              .writedata
		.pll_reconfigurar_mgmt_avalon_slave_waitrequest                      (mm_interconnect_0_pll_reconfigurar_mgmt_avalon_slave_waitrequest), //                                                              .waitrequest
		.reset_s1_address                                                    (mm_interconnect_0_reset_s1_address),                               //                                                      reset_s1.address
		.reset_s1_write                                                      (mm_interconnect_0_reset_s1_write),                                 //                                                              .write
		.reset_s1_readdata                                                   (mm_interconnect_0_reset_s1_readdata),                              //                                                              .readdata
		.reset_s1_writedata                                                  (mm_interconnect_0_reset_s1_writedata),                             //                                                              .writedata
		.reset_s1_chipselect                                                 (mm_interconnect_0_reset_s1_chipselect),                            //                                                              .chipselect
		.result0_32_bit_s1_address                                           (mm_interconnect_0_result0_32_bit_s1_address),                      //                                             result0_32_bit_s1.address
		.result0_32_bit_s1_readdata                                          (mm_interconnect_0_result0_32_bit_s1_readdata),                     //                                                              .readdata
		.result0_64_bit_down_s1_address                                      (mm_interconnect_0_result0_64_bit_down_s1_address),                 //                                        result0_64_bit_down_s1.address
		.result0_64_bit_down_s1_readdata                                     (mm_interconnect_0_result0_64_bit_down_s1_readdata),                //                                                              .readdata
		.result0_64_bit_up_s1_address                                        (mm_interconnect_0_result0_64_bit_up_s1_address),                   //                                          result0_64_bit_up_s1.address
		.result0_64_bit_up_s1_readdata                                       (mm_interconnect_0_result0_64_bit_up_s1_readdata),                  //                                                              .readdata
		.result1_32_bit_s1_address                                           (mm_interconnect_0_result1_32_bit_s1_address),                      //                                             result1_32_bit_s1.address
		.result1_32_bit_s1_readdata                                          (mm_interconnect_0_result1_32_bit_s1_readdata),                     //                                                              .readdata
		.result1_64_bit_down_s1_address                                      (mm_interconnect_0_result1_64_bit_down_s1_address),                 //                                        result1_64_bit_down_s1.address
		.result1_64_bit_down_s1_readdata                                     (mm_interconnect_0_result1_64_bit_down_s1_readdata),                //                                                              .readdata
		.result1_64_bit_up_s1_address                                        (mm_interconnect_0_result1_64_bit_up_s1_address),                   //                                          result1_64_bit_up_s1.address
		.result1_64_bit_up_s1_readdata                                       (mm_interconnect_0_result1_64_bit_up_s1_readdata)                   //                                                              .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (reset_fifos_reset),                  // reset_in1.reset
		.clk            (clk_custom_in_clk),                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_custom_in_clk),                  //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
